** Profile: "SCHEMATIC1-Buck"  [ D:\Gopal\orcad\buck-pspicefiles\schematic1\buck.sim ] 

** Creating circuit file "Buck.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../buck-pspicefiles/buck.lib" 
* From [PSPICE NETLIST] section of C:\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "C:\Cadence\SPB_16.6\tools\capture\library\MOSFET\PMOS.lib" 
.lib "C:\Cadence\SPB_16.6\tools\capture\library\MOSFET\NMOS.lib" 
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 1.5ms  0 0.53372u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
