** Profile: "SCHEMATIC1-lea"  [ f:\swati\orcad_projects\leadlag-pspicefiles\schematic1\lea.sim ] 

** Creating circuit file "lea.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Users\Rahul Bhattacharya\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 110ms 0 50us 
.MC 1000 TRAN V([VOUT]) YMAX OUTPUT ALL 
+ SAVEPARAM "F:/SIMRAN_INTERN/mcp_file/lead_1000.mcp"
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
